module cmd_fifo (
    input rstn,

    input          push_clk,
    input          io_push_valid,
    output         io_push_ready,
    input          io_push_cmd_type,
    input  [ 26:0] io_push_addr,
    input  [  5:0] io_push_burst_cnt,
    input  [127:0] io_push_wt_data,
    input  [ 15:0] io_push_wt_mask,

    input          pop_clk,
    output         io_pop_valid,
    input          io_pop_ready,
    output         io_pop_cmd_type,
    output [ 26:0] io_pop_addr,
    output [  5:0] io_pop_burst_cnt,
    output [127:0] io_pop_wt_data,
    output [ 15:0] io_pop_wt_mask
);

  // 1 + 27 + 6 + 128 + 16 = 178bits
  wire [177:0] push_data;
  wire [177:0] pop_data;

  assign push_data = {
    io_push_cmd_type, io_push_addr, io_push_burst_cnt, io_push_wt_data, io_push_wt_mask
  };
  assign {io_pop_cmd_type, io_pop_addr, io_pop_burst_cnt, io_pop_wt_data, io_pop_wt_mask} = pop_data;

  FIFO_HS_CMD fifo_hs_cmd (
      .Data (push_data),
      .Reset(~rstn),
      .WrClk(push_clk),
      .RdClk(pop_clk),
      .WrEn (io_push_valid && io_push_ready),
      .RdEn (io_pop_valid && io_pop_ready),
      .Q    (pop_data),
      .Empty(~io_push_ready),
      .Full (~io_pop_ready)
  );

endmodule
